----------------------------------------------------------------------------------
-- Company: CINVESTAV
-- Engineer: JOSE DE JESUS MORALES ROMERO
-- 
-- Create Date: 30.06.2022 11:13:14
-- Design Name: ECC163
-- Module Name: FFSquarer - Behavioral
-- Project Name: ECC163
-- Target Devices: NEXYS 4 DDR
-- Tool Versions: VIVADO 2020.2
-- Description: ELEVA AL CUADRADO UN NUMERO 
-- 
-- Dependencies: 
-- 
-- Revision: 1.0
-- Revision 0.01 - File Created
-- Additional Comments: NONE
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity FFSquarer is
    Port
    (
        -- Entradas
        A: in std_logic_vector(162 downto 0);
        -- Salidas
        C: out std_logic_vector(325 downto 0)
    );
end FFSquarer;

architecture Behavioral of FFSquarer is

begin
    C(15  downto   0) <= '0' & A(  7) & '0' & A(  6) & '0' & A(  5) & '0' & A(  4) & '0' & A(  3) & '0' &  A(  2) & '0' &  A(  1) & '0' & A(  0);
    C(31  downto  16) <= '0' & A( 15) & '0' & A( 14) & '0' & A( 13) & '0' & A( 12) & '0' & A( 11) & '0' &  A( 10) & '0' &  A(  9) & '0' & A(  8);
    C(47  downto  32) <= '0' & A( 23) & '0' & A( 22) & '0' & A( 21) & '0' & A( 20) & '0' & A( 19) & '0' &  A( 18) & '0' &  A( 17) & '0' & A( 16);
    C(63  downto  48) <= '0' & A( 31) & '0' & A( 30) & '0' & A( 29) & '0' & A( 28) & '0' & A( 27) & '0' &  A( 26) & '0' &  A( 25) & '0' & A( 24);
    C(79  downto  64) <= '0' & A( 39) & '0' & A( 38) & '0' & A( 37) & '0' & A( 36) & '0' & A( 35) & '0' &  A( 34) & '0' &  A( 33) & '0' & A( 32);
    C(95  downto  80) <= '0' & A( 47) & '0' & A( 46) & '0' & A( 45) & '0' & A( 44) & '0' & A( 43) & '0' &  A( 42) & '0' &  A( 41) & '0' & A( 40);
    C(111 downto  96) <= '0' & A( 55) & '0' & A( 54) & '0' & A( 53) & '0' & A( 52) & '0' & A( 51) & '0' &  A( 50) & '0' &  A( 49) & '0' & A( 48);
    C(127 downto 112) <= '0' & A( 63) & '0' & A( 62) & '0' & A( 61) & '0' & A( 60) & '0' & A( 59) & '0' &  A( 58) & '0' &  A( 57) & '0' & A( 56);
    C(143 downto 128) <= '0' & A( 71) & '0' & A( 70) & '0' & A( 69) & '0' & A( 68) & '0' & A( 67) & '0' &  A( 66) & '0' &  A( 65) & '0' & A( 64);
    C(159 downto 144) <= '0' & A( 79) & '0' & A( 78) & '0' & A( 77) & '0' & A( 76) & '0' & A( 75) & '0' &  A( 74) & '0' &  A( 73) & '0' & A( 72);
    C(175 downto 160) <= '0' & A( 87) & '0' & A( 86) & '0' & A( 85) & '0' & A( 84) & '0' & A( 83) & '0' &  A( 82) & '0' &  A( 81) & '0' & A( 80);
    C(191 downto 161) <= '0' & A( 95) & '0' & A( 94) & '0' & A( 93) & '0' & A( 92) & '0' & A( 91) & '0' &  A( 90) & '0' &  A( 89) & '0' & A( 88);
    C(207 downto 192) <= '0' & A(103) & '0' & A(102) & '0' & A(101) & '0' & A(100) & '0' & A( 99) & '0' &  A( 98) & '0' &  A( 97) & '0' & A( 96);
    C(223 downto 208) <= '0' & A(111) & '0' & A(110) & '0' & A(109) & '0' & A(108) & '0' & A(107) & '0' &  A(106) & '0' &  A(105) & '0' & A(104);
    C(239 downto 224) <= '0' & A(119) & '0' & A(118) & '0' & A(117) & '0' & A(116) & '0' & A(115) & '0' &  A(114) & '0' &  A(113) & '0' & A(112);
    C(255 downto 240) <= '0' & A(127) & '0' & A(126) & '0' & A(125) & '0' & A(124) & '0' & A(123) & '0' &  A(122) & '0' &  A(121) & '0' & A(120);
    C(271 downto 256) <= '0' & A(135) & '0' & A(134) & '0' & A(133) & '0' & A(132) & '0' & A(131) & '0' &  A(130) & '0' &  A(129) & '0' & A(128);
    C(287 downto 272) <= '0' & A(143) & '0' & A(142) & '0' & A(141) & '0' & A(140) & '0' & A(139) & '0' &  A(138) & '0' &  A(137) & '0' & A(136);
    C(303 downto 288) <= '0' & A(151) & '0' & A(150) & '0' & A(149) & '0' & A(148) & '0' & A(147) & '0' &  A(146) & '0' &  A(145) & '0' & A(144);
    C(319 downto 304) <= '0' & A(159) & '0' & A(158) & '0' & A(157) & '0' & A(156) & '0' & A(155) & '0' &  A(154) & '0' &  A(153) & '0' & A(152);
    C(325 downto 320) <= '0' & A(162) & '0' & A(161) & '0' & A(160);
end Behavioral;
